[aimspice]
[description]
222
Invertor 2
RC EC OUT 1K
R1 IN B 1K
Q1 OUT B 0 Tranz
.MODEL Tranz NPN TR = 5e-9 TF = 8e-9
Vin IN 0 DC 0 PULSE (0 5 0 1e-9 1e-9 1e-7 2e-7)
Vec EC 0 DC 5
Veb EB 0 DC -1
Cout OUT 0 1p
C1 IN B 50P
RB B EB 7K





[tran]
1e-9
6e-7
X
X
0
[ana]
4 2
0
1 1
1 1 -4 6
3
v(out)
v(in)
v(b)
0
1 1
1 1 -4 6
2
v(out)
v(in)
[end]
