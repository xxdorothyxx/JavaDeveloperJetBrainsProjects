[aimspice]
[description]
357
TTL-NAND

Q1A 4 3 1 Tranz
Q1B 4 3 2 Tranz
Q2 6 4 5 Tranz
Q3 7 6 8 Tranz
Q4 9 5 0 Tranz

D1 0 1 myDiode
D2 0 2 myDiode
D3 8 9 myDiode

R1 cc 3 4K
R2 cc 6 1.6K
R3 cc 7 130
R4 5 0 1K

.MODEL myDiode D TT = 5e-9
.MODEL Tranz NPN TR = 5e-9 TF = 8e-9

Vcc cc 0 DC 5 
VA 1 0 DC 5 pulse(0 5 0 1e-9 1e-9 1e-8 2e-8)
VB 2 0 DC 5

C1 9 0 15p


[dc]
1
VA
0
5
0.1
[tran]
1e-9
6e-8
X
X
0
[ana]
4 0
[end]
