[aimspice]
[description]
298
Nmos Static Invertor

m1 out in 0 0 nmos_m1 L=1u W=1u
.model nmos_m1 nmos vto = 1.5 !tensiunea de prag / tresh hold voltage

m2 d g out out nmos_m2 L=25u W=1u
.model nmos_m2 nmos vto = 2.5 !tensiunea de prag

vdd d 0 dc 5
vgg g 0 dc 7.5

vin in 0 dc 5 pulse(0 5 0 1e-10 1e-10 1e-9 2e-9) 
[dc]
1
vin
0
5
0.1
[tran]
1e-9
6e-9
X
X
0
[ana]
4 1
0
1 1
1 1 -1 6
2
v(out)
v(in)
[end]
