library ieee;
use ieee.std_logic_1164.all; 
use ieee.std_logic_unsigned.all;

entity RAM_TENTATIVA1 is
	port(A: in std_logic_vector(3 downto 0);
	CLK,CE_WR: in std_logic;
	DI: in std_logic_vector(31 downto 0);
	DO: out std_logic_vector(31 downto 0));
end RAM_TENTATIVA1; 

architecture bairam of RAM_TENTATIVA1 is
type MATRIX is array (0 to 15) of std_logic_vector(31 downto 0);
begin
	process(A,CLK,CE_WR)
	variable M: MATRIX:=("00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000010","00000000000000000000000000000011","00000000000000000000000000000100","00000000000000000000000000000101","00000000000000000000000000000110","00000000000000000000000000000111","00000000000000000000000000001000","00000000000000000000000000001001","00000000000000000000000000001010","00000000000000000000000000001011","00000000000000000000000000001100","00000000000000000000000000001101","00000000000000000000000000001110","00000000000000000000000000001111");
	begin
		if CLK'EVENT and CLK='1' then
				if CE_WR='1' then
					M(conv_integer(A)):=DI; 
				else
					DO<=M(conv_integer(A));
				end if;
		end if;
	end process;
end architecture bairam;