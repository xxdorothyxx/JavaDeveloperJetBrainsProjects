[aimspice]
[description]
152
Filter rectifier

RL 4 0 100
C1 4 0 3m
D1 1 4 Diode
D2 0 1 Diode
D3 0 3 Diode
D4 3 4 Diode

.model Diode d tt = 1e-9

Vin 1 3 sin(0 5 1k 0 0)
[tran]
1e-9
6e-3
X
X
0
[ana]
4 1
0
1 1
1 1 -1 5
3
v(4)
v(1)
v(3)
[end]
