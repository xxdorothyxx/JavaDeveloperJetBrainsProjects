[aimspice]
[description]
289
Raection regulator with no error amplifier
R1 2 Z 220
RL OUT 0 100
C1 2 0 1M
D1 1 2 DiodeS
D2 3 2 DiodeS
D3 0 3 DiodeS
D4 0 1 DiodeS
Dz 0 Z DiodeZ
Q1 2 Z OUT Tranz
.MODEL Tranz NPN TR = 1e-9 TF = 1e-9
.MODEL DiodeS D TT = 1e-9
.MODEL DiodeZ D BV = 5.6
Vin 1 3 sin(0 10 50 0 0)
[tran]
1e-9
6e-2
X
X
0
[ana]
4 1
0
1 1
1 1 -2 10
5
v(2)
v(z)
v(out)
v(1)
v(3)
[end]
