[aimspice]
[description]
94
Rectifiers
d1 1 2 myDiode
.model myDiode d tt= 1e-9
rl 2 0 100k
vin 1 0 sin ( 0 5 1k 0 0 )
[tran]
1e-9
6e-3
0
0.00001
0
[ana]
4 0
[end]
