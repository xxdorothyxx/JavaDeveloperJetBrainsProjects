[aimspice]
[description]
258
The static NOR

M1 OUT A 0 0 NMOS1 l=1u w=10u
M2 OUT B 0 0 NMOS1 l=1u w=10u
.model NMOS1 nmos vto=1.5
M3 DD GG OUT OUT NMOS2 l=10u w=1u
.model NMOS2 nmos vto=2.5

Vdd DD 0 DC 5
Vgg GG 0 DC 7.5
Va A 0 PULSE (0 5 0 1e-10 1e-10 1e-9 2e-9)
Vb B 0 DC 0
[tran]
1e-9
6e-9
X
X
0
[ana]
4 0
[end]
