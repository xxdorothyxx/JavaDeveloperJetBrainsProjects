[aimspice]
[description]
295
Reaction regulator with no error amplifier

RL 2 0 100
R1 4 5 220
C1 4 0 3m
D5 0 5 DiodeZ
D1 1 4 Diode
D2 0 1 Diode
D3 0 3 Diode
D4 3 4 Diode
Q1 4 5 2 tranzistor

.model Diode d tt = 1e-9
.model DiodeZ d bv = 6.8
.model tranzistor NPN tr = 5e-9 tf = 8e-9

Vin 1 3 sin(0 5 1k 0 0)
[end]
