[aimspice]
[description]
144
Full-wave rectifier

RL 4 0 100
D1 1 4 Diode
D2 0 1 Diode
D3 0 3 Diode
D4 3 4 Diode

.model Diode d tt = 1e-9

Vin 1 3 sin(0 5 1k 0 0)
[end]
