[aimspice]
[description]
208
Inverter with bipolar transistor

R1 IN 1 1k
C1 IN 1 15p
RB 1 EB 7k
RC EC OUT 1k
Q1 OUT 1 0 transistor

.model transistor NPN tr=5e-9 tf=8e-9
VEB EB 0 DC -1
VEC EC 0 DC 5

Vin IN 0 sin(0 5 1k 0 0)
[end]
