[aimspice]
[description]
228
Parametric regulator with Zener diode

RL 4 0 100
C1 4 0 3m
D5 0 4 DiodeZ
D1 1 4 Diode
D2 0 1 Diode
D3 0 3 Diode
D4 3 4 Diode

.model Diode d tt = 1e-9
.model DiodeZ d bv = 6.8

Vin 1 3 sin(0 5 1k 0 0)
!Vin 1 3 5

[dc]
1
Vin
0
5
0.1
[tran]
1e-9
6e-3
X
X
0
[ana]
1 1
0
1 1
1 1 -1 5
3
v(4)
v(1)
v(3)
[end]
