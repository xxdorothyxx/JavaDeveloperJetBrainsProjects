[aimspice]
[description]
215
Parametric regulator with Zenner diode
RL 2 0 100
C1 2 0 1M
D1 1 2 DiodeS
D2 3 2 DiodeS
D3 0 3 DiodeS
D4 0 1 DiodeS
Dz 0 2 DiodeZ
.MODEL DiodeS D TT = 1e-9
.MODEL DiodeZ D BV = 6.8
Vin 1 3 sin(0 10 50 0 0)
[tran]
1e-9
6e-2
X
X
0
[ana]
4 1
0
1 1
1 1 -3.44663E-29 8
1
v(2)
[end]
