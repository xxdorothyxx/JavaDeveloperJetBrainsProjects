[aimspice]
[description]
160
Rectifiers full
d1 1 2 myDiode
.model myDiode d tt= 1e-9
d2 3 2 myDiode
d3 0 3 myDiode
d4 0 1 myDiode
rl 2 0 100k
c1 2 0 0.1m
vin 1 3 sin ( 0 5 1k 0 0 )
[tran]
1e-9
6e-3
0
0.00001
0
[end]
