[aimspice]
[description]
261
NAND NMOS

M1 temp b 0 0 NMOS1 l=1u w=10u
M2 out a temp temp NMOS1 l=1u w=10u
.Model NMOS1 nmos vto=1.5

M3 dd gg out out NMOS2 l=10u w=1u
.Model NMOS2 nmos vto=2.5

Vdd dd 0 DC 5
Vgg gg 0 DC 7.5
Va a 0 pulse(0 5 0 1e-10 1e-10 1e-9 2e-9)
Vb b 0 DC 5
[tran]
1e-10
5e-9
X
X
0
[ana]
4 1
0
1 1
1 1 -1 6
3
v(b)
v(out)
v(a)
[end]
